non linearity 
.include ua741.txt 
r1 2 3 9.9776k
D1 3 4 
r2 3 1 60.4K
D2 4 1 
x1 gnd 3 5 6 4 UA741
x2 gnd 7 5 6 8 UA741
x3 gnd 9 5 6 10 UA741
x4 gnd 14 5 6 11 UA741
x5 gnd 12 5 6 2 UA741
r3 7 1 13.208k
r4 7 8 13.226k
r5 8 9 13.251k
r6 13 9 199.81k
r7 10 14 13.25k
r8 11 12 13.268k
r9 7 11 13.23k
c1 9 10 9.882n
c2 14 11 9.853n
c3 12 2 9.924n 
rv 9 10 5k
v1 5 gnd 15v
v2 6 gnd -15v
v3 13 gnd 5v
.control
tran 0.00001 0.06
plot v(2)
.endc 
.end 
