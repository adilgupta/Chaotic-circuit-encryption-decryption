non linearity 
.include ua741.txt 
r1 2 3 9.9776k
D1 3 4 
r2 3 1 60.4K
D2 4 1 
x1 gnd 3 5 6 4 UA741
x2 gnd 7 5 6 8 UA741
x3 gnd 9 5 6 10 UA741
x4 gnd 14 5 6 11 UA741
x5 gnd 12 5 6 2 UA741
r3 7 1 13.208k
r4 7 8 13.226k
r5 8 9 13.251k
r6 13 9 199.81k
r7 10 14 13.25k
r8 11 12 13.268k
r9 7 11 13.23k
c1 9 10 9.882n
c2 14 11 9.853n
c3 12 2 9.924n 
rv 9 10 20k
v1 5 gnd 20v
v2 6 gnd -15v
v3 13 gnd 5v
r10 2 15 100.31k
r11 15 16 100.06k
r12 15 17 100.12k
r13 17 18 100.31k
r14 18 19 100.24k
x6 gnd 15 5 6 17 ua741
x7 gnd 18 5 6 19 ua741
vin 16 0 sin(0 0.25 100 0 0 0)
r15 19 20 20.091k
r16 20 40 15.995k
x8 gnd 20 5 6 40 ua741
r17 50 24 9.9776k
D3 24 25 
r18 24 22 60.4K
D4 25 22 
x9 gnd 24 5 6 25 UA741
x10 gnd 28 5 6 29 UA741
x11 gnd 30 5 6 31 UA741
x12 gnd 35 5 6 32 UA741
x13 gnd 33 5 6 42 UA741
r19 28 22 13.208k
r20 28 29 13.226k
r21 29 30 13.252k
r22 34 30 199.81k
r23 31 35 13.248k
r24 32 33 13.272k
r25 28 32 13.23k
c4 30 31 9.879n
c5 35 32 9.861n
c6 33 42 9.909n 
rv2 30 31 20k
v4 34 gnd 5v
r26 42 20 80.091k
x14 gnd 41 5 6 50 ua741
r27 40 41 100k
r28 41 50 100k 
r29 17 43 100k
r30 42 43 100k
r31 43 44 100k
x15 gnd 43 5 6 44 UA741
.control
tran 0.0001 0.12
plot v(42)+V(17)
plot v(44)
.endc 
.end 
