non linearity 
.include ua741.txt 
r1 2 3 9.9776k
D1 3 4 
r2 3 1 60.4K
D2 4 1 
x1 gnd 3 5 6 4 UA741
x2 gnd 7 5 6 8 UA741
x3 gnd 9 5 6 10 UA741
x4 gnd 14 5 6 11 UA741
x5 gnd 12 5 6 2 UA741
r3 7 1 13.208k
r4 7 8 13.226k
r5 8 9 13.251k
r6 13 9 199.81k
r7 10 14 13.25k
r8 11 12 13.268k
r9 7 11 13.23k
c1 9 10 9.882n
c2 14 11 9.853n
c3 12 2 9.924n 
rv 9 10 20k
v1 5 gnd 15v
v2 6 gnd -15v
v3 13 gnd 5v
r10 2 15 100.31k
r11 15 16 100.06k
r12 15 17 100.12k
r13 17 18 100.31k
r14 18 19 100.24k
x6 gnd 15 5 6 17 ua741
x7 gnd 18 5 6 19 ua741
vin 16 0 sin(0 0.1 100 0 0 0)
.control
tran 0.0001 0.12
plot v(19)
.endc 
.end 
